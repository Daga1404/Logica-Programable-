module floor_change (
    input clk, rst, enable,
    input [4:0] selected_floor,
    output reg [0:6] HEX0, HEX1,
    output reg open_door
);
    
    
endmodule